module instruction_fetch(unextend,extended);


endmodule
